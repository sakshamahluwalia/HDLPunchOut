module enemy_meta_datapath(clock, reset_n, enable, x_pos, x_out,	y_out, c_out);
	input clock;
	input reset_n;
	input enable;
	input [7:0] x_pos;
	
	output reg [7:0] x_out;
	output reg [6:0] y_out;
	output reg c_out;
	


endmodule