module user_data(SW, clock, reset_n, block);



endmodule